// $Id: $
// File name:   tb_Arctan.sv
// Created:     4/2/2014
// Author:      Yuchen Cui
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: test bench for arctan
`timescale 1ns/1ps

module tb_Arctan();
  
  reg [15:0] x_in,y_in;
  reg [15:0] angle;
  
  Arctan DUT (
    .x_in(x_in),
    .y_in(y_in),
    .angle_out(angle)
  );
  
  initial
  begin
    #10;
    x_in = 16'b0111111111111110;
    y_in = 16'b0111111111111111;
    #200;
    x_in = 16'b0000000011111111;
    y_in = 16'b0111111110000000;
    #200;
    x_in = 16'b0100000011111111;
    y_in = 16'b0111000000000111;
    #200;
    x_in = 16'b0100000011111111;
    y_in = 16'b0111111111111111;
    #200;
    y_in = 16'b0000000011111111;
    x_in = 16'b0111110000000000;
    #200;
    y_in = 16'b0000000000000001;
    x_in = 16'b0111111111111111;
    #200;
    x_in = 16'b0000000000000011;
    y_in = 16'b0000000000000011;
    #200;
    x_in = 16'b1000000011111111;
    y_in = 16'b0111100001111111;
    #200;
    x_in = 16'b0100000011111111;
    y_in = 16'b0111111111111111;
    #200;
    x_in = 16'b0100000011111111;
    y_in = 16'b0111111111111111;
    #200;
    y_in = 16'b0000000011111111;
    x_in = 16'b0111111111111111;
    #200;
    y_in = 16'b1000000000000001;
    x_in = 16'b1111111111111111;
    #200;
    x_in = 16'b0000000000000011;
    y_in = 16'b1000000000000011;
    #200;
    x_in = 16'b0000000000000011;
    y_in = 16'b1111111111111100;
    #200;
    x_in = 16'b0000011111000011;
    y_in = 16'b1001111000000011;
    #200;
    x_in = 16'b0001111000000011;
    y_in = 16'b1000000000000011;
    #200;
    x_in = 16'b1000000000000011;
    y_in = 16'b1000000000000011;
    #200;
    x_in = 16'b1000100000000011;
    y_in = 16'b1000000000000011;
    #200;
    x_in = 16'b1000100000000011;
    y_in = 16'b1000000000000011;
  end
endmodule