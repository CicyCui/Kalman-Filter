// $Id: $
// File name:   datapath.sv
// Created:     4/15/2014
// Author:      Yuhao Chen
// Lab Section: 2
// Version:     1.0  Initial Design Entry
// Description: datapath for output
module datapath
(
  input wire [7:0] rx_write_data,
  input wire [7:0] addr,
  output reg [47:0] acc_data,
  output reg [47:0] gyro_data,
  output reg [47:0] mag_data
);





endmodule