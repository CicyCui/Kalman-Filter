// $Id: $
// File name:   tb_Preprocessor.sv
// Created:     4/9/2014
// Author:      Yuchen Cui
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: test bench for preprocessor
