// $Id: $
// File name:   Arctan.sv
// Created:     4/1/2014
// Author:      Yuchen Cui
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: arctan calculation module
module Arctan(
  input wire [15:0] x_in,
  input wire [15:0] y_in,
  output wire [15:0] angle_out
  );
  
  reg [9:0] ratio; 
  reg [15:0] x,y;
  reg [15:0] new_angle,angle,angle_complement;
  reg [15:0] num,den;
  reg [24:0] product;

  assign angle_out = new_angle;
  assign num = x < y ? x:y;
  assign den = x > y ? x:y;
  assign angle_complement =  {16'b0100000000000000} - angle; 
  assign product = 1023 * num;
  assign ratio = product / den;
  
  //output logic
  always_comb begin
    if(x_in[15] == 1'b1) begin
      x[15] = 0;
      x[14:0] = ~{x_in[14:0]} + 1'b1;
    end
  else x = x_in;
    if(y_in[15] == 1'b1) begin
      y[15] = 0;
      y[14:0] = ~{y_in[14:0]} + 1'b1;
    end
  else y = y_in;
  end
  
  
  always_comb begin
    if(x_in[14:0] == 0 )
    begin
        if(y_in[15] == 1'b0) begin //x=0 y > 0
          new_angle = 0;//0
        end
        else begin // x=0 y<0
          new_angle = {16'b1000000000000000};//180
        end
    end  
    else if ( y_in[14:0] == 0 ) begin
       if(x_in[15] == 1'b0)begin
         new_angle = {16'b0100000000000000};//90
       end
     else begin
         new_angle = {16'b1100000000000000};//270
     end
    end
    else
      begin
   if(y_in[15] == 1'b0) begin // section I and IV
      if(x_in[15] == 1'b0) begin //section I
        if( x <= y ) begin // 0-45
          new_angle = angle;
        end else begin//45 - 90
          new_angle = angle_complement;  //90-x
        end
      end else begin //section IV
        if( x <= y ) begin // 315-360
          new_angle = angle_complement + {16'b1100000000000000}; //+45*6
        end else begin //270-315
          new_angle = angle + {16'b1100000000000000}; //+45*6
        end
      end
    end else begin  //section II & III
      if(x_in[15] == 1'b0) begin //section II
        if( x <= y ) begin // 135-180
          new_angle = angle_complement + {16'b0100000000000000}; //45*2
        end else begin //90-135
          new_angle = angle + {16'b0100000000000000}; //+45*2
        end
      end else begin //section III
        if( x <= y ) begin // 180-225
          new_angle = angle + {16'b1000000000000000}; //*4
        end else begin //225-270
          new_angle = angle_complement + {16'b1000000000000000};//*4
        end
      end  
    end
  end
    
    
  end

//lookup table for arctan: precision is of step 45/1024
always_comb begin
case(ratio)  
    10'b0000000000: angle = 16'b0000000000000000;
    10'b0000000001: angle = 16'b0000000000001010;
    10'b0000000010: angle = 16'b0000000000010100;
    10'b0000000011: angle = 16'b0000000000011110;
    10'b0000000100: angle = 16'b0000000000101000;
    10'b0000000101: angle = 16'b0000000000110010;
    10'b0000000110: angle = 16'b0000000000111101;
    10'b0000000111: angle = 16'b0000000001000111;
    10'b0000001000: angle = 16'b0000000001010001;
    10'b0000001001: angle = 16'b0000000001011011;
    10'b0000001010: angle = 16'b0000000001100101;
    10'b0000001011: angle = 16'b0000000001110000;
    10'b0000001100: angle = 16'b0000000001111010;
    10'b0000001101: angle = 16'b0000000010000100;
    10'b0000001110: angle = 16'b0000000010001110;
    10'b0000001111: angle = 16'b0000000010011000;
    10'b0000010000: angle = 16'b0000000010100010;
    10'b0000010001: angle = 16'b0000000010101101;
    10'b0000010010: angle = 16'b0000000010110111;
    10'b0000010011: angle = 16'b0000000011000001;
    10'b0000010100: angle = 16'b0000000011001011;
    10'b0000010101: angle = 16'b0000000011010101;
    10'b0000010110: angle = 16'b0000000011100000;
    10'b0000010111: angle = 16'b0000000011101010;
    10'b0000011000: angle = 16'b0000000011110100;
    10'b0000011001: angle = 16'b0000000011111110;
    10'b0000011010: angle = 16'b0000000100001000;
    10'b0000011011: angle = 16'b0000000100010010;
    10'b0000011100: angle = 16'b0000000100011101;
    10'b0000011101: angle = 16'b0000000100100111;
    10'b0000011110: angle = 16'b0000000100110001;
    10'b0000011111: angle = 16'b0000000100111011;
    10'b0000100000: angle = 16'b0000000101000101;
    10'b0000100001: angle = 16'b0000000101010000;
    10'b0000100010: angle = 16'b0000000101011010;
    10'b0000100011: angle = 16'b0000000101100100;
    10'b0000100100: angle = 16'b0000000101101110;
    10'b0000100101: angle = 16'b0000000101111000;
    10'b0000100110: angle = 16'b0000000110000010;
    10'b0000100111: angle = 16'b0000000110001101;
    10'b0000101000: angle = 16'b0000000110010111;
    10'b0000101001: angle = 16'b0000000110100001;
    10'b0000101010: angle = 16'b0000000110101011;
    10'b0000101011: angle = 16'b0000000110110101;
    10'b0000101100: angle = 16'b0000000110111111;
    10'b0000101101: angle = 16'b0000000111001010;
    10'b0000101110: angle = 16'b0000000111010100;
    10'b0000101111: angle = 16'b0000000111011110;
    10'b0000110000: angle = 16'b0000000111101000;
    10'b0000110001: angle = 16'b0000000111110010;
    10'b0000110010: angle = 16'b0000000111111100;
    10'b0000110011: angle = 16'b0000001000000111;
    10'b0000110100: angle = 16'b0000001000010001;
    10'b0000110101: angle = 16'b0000001000011011;
    10'b0000110110: angle = 16'b0000001000100101;
    10'b0000110111: angle = 16'b0000001000101111;
    10'b0000111000: angle = 16'b0000001000111001;
    10'b0000111001: angle = 16'b0000001001000011;
    10'b0000111010: angle = 16'b0000001001001110;
    10'b0000111011: angle = 16'b0000001001011000;
    10'b0000111100: angle = 16'b0000001001100010;
    10'b0000111101: angle = 16'b0000001001101100;
    10'b0000111110: angle = 16'b0000001001110110;
    10'b0000111111: angle = 16'b0000001010000000;
    10'b0001000000: angle = 16'b0000001010001011;
    10'b0001000001: angle = 16'b0000001010010101;
    10'b0001000010: angle = 16'b0000001010011111;
    10'b0001000011: angle = 16'b0000001010101001;
    10'b0001000100: angle = 16'b0000001010110011;
    10'b0001000101: angle = 16'b0000001010111101;
    10'b0001000110: angle = 16'b0000001011000111;
    10'b0001000111: angle = 16'b0000001011010010;
    10'b0001001000: angle = 16'b0000001011011100;
    10'b0001001001: angle = 16'b0000001011100110;
    10'b0001001010: angle = 16'b0000001011110000;
    10'b0001001011: angle = 16'b0000001011111010;
    10'b0001001100: angle = 16'b0000001100000100;
    10'b0001001101: angle = 16'b0000001100001110;
    10'b0001001110: angle = 16'b0000001100011000;
    10'b0001001111: angle = 16'b0000001100100011;
    10'b0001010000: angle = 16'b0000001100101101;
    10'b0001010001: angle = 16'b0000001100110111;
    10'b0001010010: angle = 16'b0000001101000001;
    10'b0001010011: angle = 16'b0000001101001011;
    10'b0001010100: angle = 16'b0000001101010101;
    10'b0001010101: angle = 16'b0000001101011111;
    10'b0001010110: angle = 16'b0000001101101001;
    10'b0001010111: angle = 16'b0000001101110100;
    10'b0001011000: angle = 16'b0000001101111110;
    10'b0001011001: angle = 16'b0000001110001000;
    10'b0001011010: angle = 16'b0000001110010010;
    10'b0001011011: angle = 16'b0000001110011100;
    10'b0001011100: angle = 16'b0000001110100110;
    10'b0001011101: angle = 16'b0000001110110000;
    10'b0001011110: angle = 16'b0000001110111010;
    10'b0001011111: angle = 16'b0000001111000100;
    10'b0001100000: angle = 16'b0000001111001110;
    10'b0001100001: angle = 16'b0000001111011001;
    10'b0001100010: angle = 16'b0000001111100011;
    10'b0001100011: angle = 16'b0000001111101101;
    10'b0001100100: angle = 16'b0000001111110111;
    10'b0001100101: angle = 16'b0000010000000001;
    10'b0001100110: angle = 16'b0000010000001011;
    10'b0001100111: angle = 16'b0000010000010101;
    10'b0001101000: angle = 16'b0000010000011111;
    10'b0001101001: angle = 16'b0000010000101001;
    10'b0001101010: angle = 16'b0000010000110011;
    10'b0001101011: angle = 16'b0000010000111101;
    10'b0001101100: angle = 16'b0000010001001000;
    10'b0001101101: angle = 16'b0000010001010010;
    10'b0001101110: angle = 16'b0000010001011100;
    10'b0001101111: angle = 16'b0000010001100110;
    10'b0001110000: angle = 16'b0000010001110000;
    10'b0001110001: angle = 16'b0000010001111010;
    10'b0001110010: angle = 16'b0000010010000100;
    10'b0001110011: angle = 16'b0000010010001110;
    10'b0001110100: angle = 16'b0000010010011000;
    10'b0001110101: angle = 16'b0000010010100010;
    10'b0001110110: angle = 16'b0000010010101100;
    10'b0001110111: angle = 16'b0000010010110110;
    10'b0001111000: angle = 16'b0000010011000000;
    10'b0001111001: angle = 16'b0000010011001010;
    10'b0001111010: angle = 16'b0000010011010100;
    10'b0001111011: angle = 16'b0000010011011110;
    10'b0001111100: angle = 16'b0000010011101000;
    10'b0001111101: angle = 16'b0000010011110010;
    10'b0001111110: angle = 16'b0000010011111101;
    10'b0001111111: angle = 16'b0000010100000111;
    10'b0010000000: angle = 16'b0000010100010001;
    10'b0010000001: angle = 16'b0000010100011011;
    10'b0010000010: angle = 16'b0000010100100101;
    10'b0010000011: angle = 16'b0000010100101111;
    10'b0010000100: angle = 16'b0000010100111001;
    10'b0010000101: angle = 16'b0000010101000011;
    10'b0010000110: angle = 16'b0000010101001101;
    10'b0010000111: angle = 16'b0000010101010111;
    10'b0010001000: angle = 16'b0000010101100001;
    10'b0010001001: angle = 16'b0000010101101011;
    10'b0010001010: angle = 16'b0000010101110101;
    10'b0010001011: angle = 16'b0000010101111111;
    10'b0010001100: angle = 16'b0000010110001001;
    10'b0010001101: angle = 16'b0000010110010011;
    10'b0010001110: angle = 16'b0000010110011101;
    10'b0010001111: angle = 16'b0000010110100111;
    10'b0010010000: angle = 16'b0000010110110001;
    10'b0010010001: angle = 16'b0000010110111011;
    10'b0010010010: angle = 16'b0000010111000101;
    10'b0010010011: angle = 16'b0000010111001111;
    10'b0010010100: angle = 16'b0000010111011001;
    10'b0010010101: angle = 16'b0000010111100011;
    10'b0010010110: angle = 16'b0000010111101101;
    10'b0010010111: angle = 16'b0000010111110111;
    10'b0010011000: angle = 16'b0000011000000001;
    10'b0010011001: angle = 16'b0000011000001011;
    10'b0010011010: angle = 16'b0000011000010100;
    10'b0010011011: angle = 16'b0000011000011110;
    10'b0010011100: angle = 16'b0000011000101000;
    10'b0010011101: angle = 16'b0000011000110010;
    10'b0010011110: angle = 16'b0000011000111100;
    10'b0010011111: angle = 16'b0000011001000110;
    10'b0010100000: angle = 16'b0000011001010000;
    10'b0010100001: angle = 16'b0000011001011010;
    10'b0010100010: angle = 16'b0000011001100100;
    10'b0010100011: angle = 16'b0000011001101110;
    10'b0010100100: angle = 16'b0000011001111000;
    10'b0010100101: angle = 16'b0000011010000010;
    10'b0010100110: angle = 16'b0000011010001100;
    10'b0010100111: angle = 16'b0000011010010110;
    10'b0010101000: angle = 16'b0000011010100000;
    10'b0010101001: angle = 16'b0000011010101010;
    10'b0010101010: angle = 16'b0000011010110011;
    10'b0010101011: angle = 16'b0000011010111101;
    10'b0010101100: angle = 16'b0000011011000111;
    10'b0010101101: angle = 16'b0000011011010001;
    10'b0010101110: angle = 16'b0000011011011011;
    10'b0010101111: angle = 16'b0000011011100101;
    10'b0010110000: angle = 16'b0000011011101111;
    10'b0010110001: angle = 16'b0000011011111001;
    10'b0010110010: angle = 16'b0000011100000011;
    10'b0010110011: angle = 16'b0000011100001101;
    10'b0010110100: angle = 16'b0000011100010110;
    10'b0010110101: angle = 16'b0000011100100000;
    10'b0010110110: angle = 16'b0000011100101010;
    10'b0010110111: angle = 16'b0000011100110100;
    10'b0010111000: angle = 16'b0000011100111110;
    10'b0010111001: angle = 16'b0000011101001000;
    10'b0010111010: angle = 16'b0000011101010010;
    10'b0010111011: angle = 16'b0000011101011100;
    10'b0010111100: angle = 16'b0000011101100101;
    10'b0010111101: angle = 16'b0000011101101111;
    10'b0010111110: angle = 16'b0000011101111001;
    10'b0010111111: angle = 16'b0000011110000011;
    10'b0011000000: angle = 16'b0000011110001101;
    10'b0011000001: angle = 16'b0000011110010111;
    10'b0011000010: angle = 16'b0000011110100000;
    10'b0011000011: angle = 16'b0000011110101010;
    10'b0011000100: angle = 16'b0000011110110100;
    10'b0011000101: angle = 16'b0000011110111110;
    10'b0011000110: angle = 16'b0000011111001000;
    10'b0011000111: angle = 16'b0000011111010010;
    10'b0011001000: angle = 16'b0000011111011011;
    10'b0011001001: angle = 16'b0000011111100101;
    10'b0011001010: angle = 16'b0000011111101111;
    10'b0011001011: angle = 16'b0000011111111001;
    10'b0011001100: angle = 16'b0000100000000011;
    10'b0011001101: angle = 16'b0000100000001100;
    10'b0011001110: angle = 16'b0000100000010110;
    10'b0011001111: angle = 16'b0000100000100000;
    10'b0011010000: angle = 16'b0000100000101010;
    10'b0011010001: angle = 16'b0000100000110100;
    10'b0011010010: angle = 16'b0000100000111101;
    10'b0011010011: angle = 16'b0000100001000111;
    10'b0011010100: angle = 16'b0000100001010001;
    10'b0011010101: angle = 16'b0000100001011011;
    10'b0011010110: angle = 16'b0000100001100100;
    10'b0011010111: angle = 16'b0000100001101110;
    10'b0011011000: angle = 16'b0000100001111000;
    10'b0011011001: angle = 16'b0000100010000010;
    10'b0011011010: angle = 16'b0000100010001011;
    10'b0011011011: angle = 16'b0000100010010101;
    10'b0011011100: angle = 16'b0000100010011111;
    10'b0011011101: angle = 16'b0000100010101001;
    10'b0011011110: angle = 16'b0000100010110010;
    10'b0011011111: angle = 16'b0000100010111100;
    10'b0011100000: angle = 16'b0000100011000110;
    10'b0011100001: angle = 16'b0000100011001111;
    10'b0011100010: angle = 16'b0000100011011001;
    10'b0011100011: angle = 16'b0000100011100011;
    10'b0011100100: angle = 16'b0000100011101101;
    10'b0011100101: angle = 16'b0000100011110110;
    10'b0011100110: angle = 16'b0000100100000000;
    10'b0011100111: angle = 16'b0000100100001010;
    10'b0011101000: angle = 16'b0000100100010011;
    10'b0011101001: angle = 16'b0000100100011101;
    10'b0011101010: angle = 16'b0000100100100111;
    10'b0011101011: angle = 16'b0000100100110000;
    10'b0011101100: angle = 16'b0000100100111010;
    10'b0011101101: angle = 16'b0000100101000100;
    10'b0011101110: angle = 16'b0000100101001101;
    10'b0011101111: angle = 16'b0000100101010111;
    10'b0011110000: angle = 16'b0000100101100001;
    10'b0011110001: angle = 16'b0000100101101010;
    10'b0011110010: angle = 16'b0000100101110100;
    10'b0011110011: angle = 16'b0000100101111110;
    10'b0011110100: angle = 16'b0000100110000111;
    10'b0011110101: angle = 16'b0000100110010001;
    10'b0011110110: angle = 16'b0000100110011011;
    10'b0011110111: angle = 16'b0000100110100100;
    10'b0011111000: angle = 16'b0000100110101110;
    10'b0011111001: angle = 16'b0000100110111000;
    10'b0011111010: angle = 16'b0000100111000001;
    10'b0011111011: angle = 16'b0000100111001011;
    10'b0011111100: angle = 16'b0000100111010100;
    10'b0011111101: angle = 16'b0000100111011110;
    10'b0011111110: angle = 16'b0000100111101000;
    10'b0011111111: angle = 16'b0000100111110001;
    10'b0100000000: angle = 16'b0000100111111011;
    10'b0100000001: angle = 16'b0000101000000100;
    10'b0100000010: angle = 16'b0000101000001110;
    10'b0100000011: angle = 16'b0000101000010111;
    10'b0100000100: angle = 16'b0000101000100001;
    10'b0100000101: angle = 16'b0000101000101011;
    10'b0100000110: angle = 16'b0000101000110100;
    10'b0100000111: angle = 16'b0000101000111110;
    10'b0100001000: angle = 16'b0000101001000111;
    10'b0100001001: angle = 16'b0000101001010001;
    10'b0100001010: angle = 16'b0000101001011010;
    10'b0100001011: angle = 16'b0000101001100100;
    10'b0100001100: angle = 16'b0000101001101101;
    10'b0100001101: angle = 16'b0000101001110111;
    10'b0100001110: angle = 16'b0000101010000000;
    10'b0100001111: angle = 16'b0000101010001010;
    10'b0100010000: angle = 16'b0000101010010100;
    10'b0100010001: angle = 16'b0000101010011101;
    10'b0100010010: angle = 16'b0000101010100111;
    10'b0100010011: angle = 16'b0000101010110000;
    10'b0100010100: angle = 16'b0000101010111010;
    10'b0100010101: angle = 16'b0000101011000011;
    10'b0100010110: angle = 16'b0000101011001101;
    10'b0100010111: angle = 16'b0000101011010110;
    10'b0100011000: angle = 16'b0000101011100000;
    10'b0100011001: angle = 16'b0000101011101001;
    10'b0100011010: angle = 16'b0000101011110010;
    10'b0100011011: angle = 16'b0000101011111100;
    10'b0100011100: angle = 16'b0000101100000101;
    10'b0100011101: angle = 16'b0000101100001111;
    10'b0100011110: angle = 16'b0000101100011000;
    10'b0100011111: angle = 16'b0000101100100010;
    10'b0100100000: angle = 16'b0000101100101011;
    10'b0100100001: angle = 16'b0000101100110101;
    10'b0100100010: angle = 16'b0000101100111110;
    10'b0100100011: angle = 16'b0000101101000111;
    10'b0100100100: angle = 16'b0000101101010001;
    10'b0100100101: angle = 16'b0000101101011010;
    10'b0100100110: angle = 16'b0000101101100100;
    10'b0100100111: angle = 16'b0000101101101101;
    10'b0100101000: angle = 16'b0000101101110111;
    10'b0100101001: angle = 16'b0000101110000000;
    10'b0100101010: angle = 16'b0000101110001001;
    10'b0100101011: angle = 16'b0000101110010011;
    10'b0100101100: angle = 16'b0000101110011100;
    10'b0100101101: angle = 16'b0000101110100101;
    10'b0100101110: angle = 16'b0000101110101111;
    10'b0100101111: angle = 16'b0000101110111000;
    10'b0100110000: angle = 16'b0000101111000010;
    10'b0100110001: angle = 16'b0000101111001011;
    10'b0100110010: angle = 16'b0000101111010100;
    10'b0100110011: angle = 16'b0000101111011110;
    10'b0100110100: angle = 16'b0000101111100111;
    10'b0100110101: angle = 16'b0000101111110000;
    10'b0100110110: angle = 16'b0000101111111010;
    10'b0100110111: angle = 16'b0000110000000011;
    10'b0100111000: angle = 16'b0000110000001100;
    10'b0100111001: angle = 16'b0000110000010110;
    10'b0100111010: angle = 16'b0000110000011111;
    10'b0100111011: angle = 16'b0000110000101000;
    10'b0100111100: angle = 16'b0000110000110010;
    10'b0100111101: angle = 16'b0000110000111011;
    10'b0100111110: angle = 16'b0000110001000100;
    10'b0100111111: angle = 16'b0000110001001101;
    10'b0101000000: angle = 16'b0000110001010111;
    10'b0101000001: angle = 16'b0000110001100000;
    10'b0101000010: angle = 16'b0000110001101001;
    10'b0101000011: angle = 16'b0000110001110011;
    10'b0101000100: angle = 16'b0000110001111100;
    10'b0101000101: angle = 16'b0000110010000101;
    10'b0101000110: angle = 16'b0000110010001110;
    10'b0101000111: angle = 16'b0000110010011000;
    10'b0101001000: angle = 16'b0000110010100001;
    10'b0101001001: angle = 16'b0000110010101010;
    10'b0101001010: angle = 16'b0000110010110011;
    10'b0101001011: angle = 16'b0000110010111100;
    10'b0101001100: angle = 16'b0000110011000110;
    10'b0101001101: angle = 16'b0000110011001111;
    10'b0101001110: angle = 16'b0000110011011000;
    10'b0101001111: angle = 16'b0000110011100001;
    10'b0101010000: angle = 16'b0000110011101011;
    10'b0101010001: angle = 16'b0000110011110100;
    10'b0101010010: angle = 16'b0000110011111101;
    10'b0101010011: angle = 16'b0000110100000110;
    10'b0101010100: angle = 16'b0000110100001111;
    10'b0101010101: angle = 16'b0000110100011000;
    10'b0101010110: angle = 16'b0000110100100010;
    10'b0101010111: angle = 16'b0000110100101011;
    10'b0101011000: angle = 16'b0000110100110100;
    10'b0101011001: angle = 16'b0000110100111101;
    10'b0101011010: angle = 16'b0000110101000110;
    10'b0101011011: angle = 16'b0000110101001111;
    10'b0101011100: angle = 16'b0000110101011000;
    10'b0101011101: angle = 16'b0000110101100010;
    10'b0101011110: angle = 16'b0000110101101011;
    10'b0101011111: angle = 16'b0000110101110100;
    10'b0101100000: angle = 16'b0000110101111101;
    10'b0101100001: angle = 16'b0000110110000110;
    10'b0101100010: angle = 16'b0000110110001111;
    10'b0101100011: angle = 16'b0000110110011000;
    10'b0101100100: angle = 16'b0000110110100001;
    10'b0101100101: angle = 16'b0000110110101010;
    10'b0101100110: angle = 16'b0000110110110100;
    10'b0101100111: angle = 16'b0000110110111101;
    10'b0101101000: angle = 16'b0000110111000110;
    10'b0101101001: angle = 16'b0000110111001111;
    10'b0101101010: angle = 16'b0000110111011000;
    10'b0101101011: angle = 16'b0000110111100001;
    10'b0101101100: angle = 16'b0000110111101010;
    10'b0101101101: angle = 16'b0000110111110011;
    10'b0101101110: angle = 16'b0000110111111100;
    10'b0101101111: angle = 16'b0000111000000101;
    10'b0101110000: angle = 16'b0000111000001110;
    10'b0101110001: angle = 16'b0000111000010111;
    10'b0101110010: angle = 16'b0000111000100000;
    10'b0101110011: angle = 16'b0000111000101001;
    10'b0101110100: angle = 16'b0000111000110010;
    10'b0101110101: angle = 16'b0000111000111011;
    10'b0101110110: angle = 16'b0000111001000100;
    10'b0101110111: angle = 16'b0000111001001101;
    10'b0101111000: angle = 16'b0000111001010110;
    10'b0101111001: angle = 16'b0000111001011111;
    10'b0101111010: angle = 16'b0000111001101000;
    10'b0101111011: angle = 16'b0000111001110001;
    10'b0101111100: angle = 16'b0000111001111010;
    10'b0101111101: angle = 16'b0000111010000011;
    10'b0101111110: angle = 16'b0000111010001100;
    10'b0101111111: angle = 16'b0000111010010101;
    10'b0110000000: angle = 16'b0000111010011110;
    10'b0110000001: angle = 16'b0000111010100111;
    10'b0110000010: angle = 16'b0000111010101111;
    10'b0110000011: angle = 16'b0000111010111000;
    10'b0110000100: angle = 16'b0000111011000001;
    10'b0110000101: angle = 16'b0000111011001010;
    10'b0110000110: angle = 16'b0000111011010011;
    10'b0110000111: angle = 16'b0000111011011100;
    10'b0110001000: angle = 16'b0000111011100101;
    10'b0110001001: angle = 16'b0000111011101110;
    10'b0110001010: angle = 16'b0000111011110111;
    10'b0110001011: angle = 16'b0000111011111111;
    10'b0110001100: angle = 16'b0000111100001000;
    10'b0110001101: angle = 16'b0000111100010001;
    10'b0110001110: angle = 16'b0000111100011010;
    10'b0110001111: angle = 16'b0000111100100011;
    10'b0110010000: angle = 16'b0000111100101100;
    10'b0110010001: angle = 16'b0000111100110101;
    10'b0110010010: angle = 16'b0000111100111101;
    10'b0110010011: angle = 16'b0000111101000110;
    10'b0110010100: angle = 16'b0000111101001111;
    10'b0110010101: angle = 16'b0000111101011000;
    10'b0110010110: angle = 16'b0000111101100001;
    10'b0110010111: angle = 16'b0000111101101001;
    10'b0110011000: angle = 16'b0000111101110010;
    10'b0110011001: angle = 16'b0000111101111011;
    10'b0110011010: angle = 16'b0000111110000100;
    10'b0110011011: angle = 16'b0000111110001101;
    10'b0110011100: angle = 16'b0000111110010101;
    10'b0110011101: angle = 16'b0000111110011110;
    10'b0110011110: angle = 16'b0000111110100111;
    10'b0110011111: angle = 16'b0000111110110000;
    10'b0110100000: angle = 16'b0000111110111000;
    10'b0110100001: angle = 16'b0000111111000001;
    10'b0110100010: angle = 16'b0000111111001010;
    10'b0110100011: angle = 16'b0000111111010011;
    10'b0110100100: angle = 16'b0000111111011011;
    10'b0110100101: angle = 16'b0000111111100100;
    10'b0110100110: angle = 16'b0000111111101101;
    10'b0110100111: angle = 16'b0000111111110101;
    10'b0110101000: angle = 16'b0000111111111110;
    10'b0110101001: angle = 16'b0001000000000111;
    10'b0110101010: angle = 16'b0001000000010000;
    10'b0110101011: angle = 16'b0001000000011000;
    10'b0110101100: angle = 16'b0001000000100001;
    10'b0110101101: angle = 16'b0001000000101010;
    10'b0110101110: angle = 16'b0001000000110010;
    10'b0110101111: angle = 16'b0001000000111011;
    10'b0110110000: angle = 16'b0001000001000100;
    10'b0110110001: angle = 16'b0001000001001100;
    10'b0110110010: angle = 16'b0001000001010101;
    10'b0110110011: angle = 16'b0001000001011101;
    10'b0110110100: angle = 16'b0001000001100110;
    10'b0110110101: angle = 16'b0001000001101111;
    10'b0110110110: angle = 16'b0001000001110111;
    10'b0110110111: angle = 16'b0001000010000000;
    10'b0110111000: angle = 16'b0001000010001001;
    10'b0110111001: angle = 16'b0001000010010001;
    10'b0110111010: angle = 16'b0001000010011010;
    10'b0110111011: angle = 16'b0001000010100010;
    10'b0110111100: angle = 16'b0001000010101011;
    10'b0110111101: angle = 16'b0001000010110011;
    10'b0110111110: angle = 16'b0001000010111100;
    10'b0110111111: angle = 16'b0001000011000101;
    10'b0111000000: angle = 16'b0001000011001101;
    10'b0111000001: angle = 16'b0001000011010110;
    10'b0111000010: angle = 16'b0001000011011110;
    10'b0111000011: angle = 16'b0001000011100111;
    10'b0111000100: angle = 16'b0001000011101111;
    10'b0111000101: angle = 16'b0001000011111000;
    10'b0111000110: angle = 16'b0001000100000000;
    10'b0111000111: angle = 16'b0001000100001001;
    10'b0111001000: angle = 16'b0001000100010001;
    10'b0111001001: angle = 16'b0001000100011010;
    10'b0111001010: angle = 16'b0001000100100010;
    10'b0111001011: angle = 16'b0001000100101011;
    10'b0111001100: angle = 16'b0001000100110011;
    10'b0111001101: angle = 16'b0001000100111100;
    10'b0111001110: angle = 16'b0001000101000100;
    10'b0111001111: angle = 16'b0001000101001101;
    10'b0111010000: angle = 16'b0001000101010101;
    10'b0111010001: angle = 16'b0001000101011110;
    10'b0111010010: angle = 16'b0001000101100110;
    10'b0111010011: angle = 16'b0001000101101110;
    10'b0111010100: angle = 16'b0001000101110111;
    10'b0111010101: angle = 16'b0001000101111111;
    10'b0111010110: angle = 16'b0001000110001000;
    10'b0111010111: angle = 16'b0001000110010000;
    10'b0111011000: angle = 16'b0001000110011001;
    10'b0111011001: angle = 16'b0001000110100001;
    10'b0111011010: angle = 16'b0001000110101001;
    10'b0111011011: angle = 16'b0001000110110010;
    10'b0111011100: angle = 16'b0001000110111010;
    10'b0111011101: angle = 16'b0001000111000010;
    10'b0111011110: angle = 16'b0001000111001011;
    10'b0111011111: angle = 16'b0001000111010011;
    10'b0111100000: angle = 16'b0001000111011100;
    10'b0111100001: angle = 16'b0001000111100100;
    10'b0111100010: angle = 16'b0001000111101100;
    10'b0111100011: angle = 16'b0001000111110101;
    10'b0111100100: angle = 16'b0001000111111101;
    10'b0111100101: angle = 16'b0001001000000101;
    10'b0111100110: angle = 16'b0001001000001110;
    10'b0111100111: angle = 16'b0001001000010110;
    10'b0111101000: angle = 16'b0001001000011110;
    10'b0111101001: angle = 16'b0001001000100110;
    10'b0111101010: angle = 16'b0001001000101111;
    10'b0111101011: angle = 16'b0001001000110111;
    10'b0111101100: angle = 16'b0001001000111111;
    10'b0111101101: angle = 16'b0001001001001000;
    10'b0111101110: angle = 16'b0001001001010000;
    10'b0111101111: angle = 16'b0001001001011000;
    10'b0111110000: angle = 16'b0001001001100000;
    10'b0111110001: angle = 16'b0001001001101001;
    10'b0111110010: angle = 16'b0001001001110001;
    10'b0111110011: angle = 16'b0001001001111001;
    10'b0111110100: angle = 16'b0001001010000001;
    10'b0111110101: angle = 16'b0001001010001001;
    10'b0111110110: angle = 16'b0001001010010010;
    10'b0111110111: angle = 16'b0001001010011010;
    10'b0111111000: angle = 16'b0001001010100010;
    10'b0111111001: angle = 16'b0001001010101010;
    10'b0111111010: angle = 16'b0001001010110011;
    10'b0111111011: angle = 16'b0001001010111011;
    10'b0111111100: angle = 16'b0001001011000011;
    10'b0111111101: angle = 16'b0001001011001011;
    10'b0111111110: angle = 16'b0001001011010011;
    10'b0111111111: angle = 16'b0001001011011011;
    10'b1000000000: angle = 16'b0001001011100100;
    10'b1000000001: angle = 16'b0001001011101100;
    10'b1000000010: angle = 16'b0001001011110100;
    10'b1000000011: angle = 16'b0001001011111100;
    10'b1000000100: angle = 16'b0001001100000100;
    10'b1000000101: angle = 16'b0001001100001100;
    10'b1000000110: angle = 16'b0001001100010100;
    10'b1000000111: angle = 16'b0001001100011100;
    10'b1000001000: angle = 16'b0001001100100101;
    10'b1000001001: angle = 16'b0001001100101101;
    10'b1000001010: angle = 16'b0001001100110101;
    10'b1000001011: angle = 16'b0001001100111101;
    10'b1000001100: angle = 16'b0001001101000101;
    10'b1000001101: angle = 16'b0001001101001101;
    10'b1000001110: angle = 16'b0001001101010101;
    10'b1000001111: angle = 16'b0001001101011101;
    10'b1000010000: angle = 16'b0001001101100101;
    10'b1000010001: angle = 16'b0001001101101101;
    10'b1000010010: angle = 16'b0001001101110101;
    10'b1000010011: angle = 16'b0001001101111101;
    10'b1000010100: angle = 16'b0001001110000101;
    10'b1000010101: angle = 16'b0001001110001101;
    10'b1000010110: angle = 16'b0001001110010101;
    10'b1000010111: angle = 16'b0001001110011101;
    10'b1000011000: angle = 16'b0001001110100101;
    10'b1000011001: angle = 16'b0001001110101101;
    10'b1000011010: angle = 16'b0001001110110101;
    10'b1000011011: angle = 16'b0001001110111101;
    10'b1000011100: angle = 16'b0001001111000101;
    10'b1000011101: angle = 16'b0001001111001101;
    10'b1000011110: angle = 16'b0001001111010101;
    10'b1000011111: angle = 16'b0001001111011101;
    10'b1000100000: angle = 16'b0001001111100101;
    10'b1000100001: angle = 16'b0001001111101101;
    10'b1000100010: angle = 16'b0001001111110101;
    10'b1000100011: angle = 16'b0001001111111101;
    10'b1000100100: angle = 16'b0001010000000101;
    10'b1000100101: angle = 16'b0001010000001101;
    10'b1000100110: angle = 16'b0001010000010101;
    10'b1000100111: angle = 16'b0001010000011100;
    10'b1000101000: angle = 16'b0001010000100100;
    10'b1000101001: angle = 16'b0001010000101100;
    10'b1000101010: angle = 16'b0001010000110100;
    10'b1000101011: angle = 16'b0001010000111100;
    10'b1000101100: angle = 16'b0001010001000100;
    10'b1000101101: angle = 16'b0001010001001100;
    10'b1000101110: angle = 16'b0001010001010100;
    10'b1000101111: angle = 16'b0001010001011011;
    10'b1000110000: angle = 16'b0001010001100011;
    10'b1000110001: angle = 16'b0001010001101011;
    10'b1000110010: angle = 16'b0001010001110011;
    10'b1000110011: angle = 16'b0001010001111011;
    10'b1000110100: angle = 16'b0001010010000011;
    10'b1000110101: angle = 16'b0001010010001010;
    10'b1000110110: angle = 16'b0001010010010010;
    10'b1000110111: angle = 16'b0001010010011010;
    10'b1000111000: angle = 16'b0001010010100010;
    10'b1000111001: angle = 16'b0001010010101010;
    10'b1000111010: angle = 16'b0001010010110001;
    10'b1000111011: angle = 16'b0001010010111001;
    10'b1000111100: angle = 16'b0001010011000001;
    10'b1000111101: angle = 16'b0001010011001001;
    10'b1000111110: angle = 16'b0001010011010000;
    10'b1000111111: angle = 16'b0001010011011000;
    10'b1001000000: angle = 16'b0001010011100000;
    10'b1001000001: angle = 16'b0001010011101000;
    10'b1001000010: angle = 16'b0001010011101111;
    10'b1001000011: angle = 16'b0001010011110111;
    10'b1001000100: angle = 16'b0001010011111111;
    10'b1001000101: angle = 16'b0001010100000111;
    10'b1001000110: angle = 16'b0001010100001110;
    10'b1001000111: angle = 16'b0001010100010110;
    10'b1001001000: angle = 16'b0001010100011110;
    10'b1001001001: angle = 16'b0001010100100101;
    10'b1001001010: angle = 16'b0001010100101101;
    10'b1001001011: angle = 16'b0001010100110101;
    10'b1001001100: angle = 16'b0001010100111100;
    10'b1001001101: angle = 16'b0001010101000100;
    10'b1001001110: angle = 16'b0001010101001100;
    10'b1001001111: angle = 16'b0001010101010011;
    10'b1001010000: angle = 16'b0001010101011011;
    10'b1001010001: angle = 16'b0001010101100011;
    10'b1001010010: angle = 16'b0001010101101010;
    10'b1001010011: angle = 16'b0001010101110010;
    10'b1001010100: angle = 16'b0001010101111001;
    10'b1001010101: angle = 16'b0001010110000001;
    10'b1001010110: angle = 16'b0001010110001001;
    10'b1001010111: angle = 16'b0001010110010000;
    10'b1001011000: angle = 16'b0001010110011000;
    10'b1001011001: angle = 16'b0001010110011111;
    10'b1001011010: angle = 16'b0001010110100111;
    10'b1001011011: angle = 16'b0001010110101110;
    10'b1001011100: angle = 16'b0001010110110110;
    10'b1001011101: angle = 16'b0001010110111110;
    10'b1001011110: angle = 16'b0001010111000101;
    10'b1001011111: angle = 16'b0001010111001101;
    10'b1001100000: angle = 16'b0001010111010100;
    10'b1001100001: angle = 16'b0001010111011100;
    10'b1001100010: angle = 16'b0001010111100011;
    10'b1001100011: angle = 16'b0001010111101011;
    10'b1001100100: angle = 16'b0001010111110010;
    10'b1001100101: angle = 16'b0001010111111010;
    10'b1001100110: angle = 16'b0001011000000001;
    10'b1001100111: angle = 16'b0001011000001001;
    10'b1001101000: angle = 16'b0001011000010000;
    10'b1001101001: angle = 16'b0001011000011000;
    10'b1001101010: angle = 16'b0001011000011111;
    10'b1001101011: angle = 16'b0001011000100111;
    10'b1001101100: angle = 16'b0001011000101110;
    10'b1001101101: angle = 16'b0001011000110110;
    10'b1001101110: angle = 16'b0001011000111101;
    10'b1001101111: angle = 16'b0001011001000100;
    10'b1001110000: angle = 16'b0001011001001100;
    10'b1001110001: angle = 16'b0001011001010011;
    10'b1001110010: angle = 16'b0001011001011011;
    10'b1001110011: angle = 16'b0001011001100010;
    10'b1001110100: angle = 16'b0001011001101010;
    10'b1001110101: angle = 16'b0001011001110001;
    10'b1001110110: angle = 16'b0001011001111000;
    10'b1001110111: angle = 16'b0001011010000000;
    10'b1001111000: angle = 16'b0001011010000111;
    10'b1001111001: angle = 16'b0001011010001110;
    10'b1001111010: angle = 16'b0001011010010110;
    10'b1001111011: angle = 16'b0001011010011101;
    10'b1001111100: angle = 16'b0001011010100101;
    10'b1001111101: angle = 16'b0001011010101100;
    10'b1001111110: angle = 16'b0001011010110011;
    10'b1001111111: angle = 16'b0001011010111011;
    10'b1010000000: angle = 16'b0001011011000010;
    10'b1010000001: angle = 16'b0001011011001001;
    10'b1010000010: angle = 16'b0001011011010001;
    10'b1010000011: angle = 16'b0001011011011000;
    10'b1010000100: angle = 16'b0001011011011111;
    10'b1010000101: angle = 16'b0001011011100110;
    10'b1010000110: angle = 16'b0001011011101110;
    10'b1010000111: angle = 16'b0001011011110101;
    10'b1010001000: angle = 16'b0001011011111100;
    10'b1010001001: angle = 16'b0001011100000100;
    10'b1010001010: angle = 16'b0001011100001011;
    10'b1010001011: angle = 16'b0001011100010010;
    10'b1010001100: angle = 16'b0001011100011001;
    10'b1010001101: angle = 16'b0001011100100001;
    10'b1010001110: angle = 16'b0001011100101000;
    10'b1010001111: angle = 16'b0001011100101111;
    10'b1010010000: angle = 16'b0001011100110110;
    10'b1010010001: angle = 16'b0001011100111101;
    10'b1010010010: angle = 16'b0001011101000101;
    10'b1010010011: angle = 16'b0001011101001100;
    10'b1010010100: angle = 16'b0001011101010011;
    10'b1010010101: angle = 16'b0001011101011010;
    10'b1010010110: angle = 16'b0001011101100001;
    10'b1010010111: angle = 16'b0001011101101001;
    10'b1010011000: angle = 16'b0001011101110000;
    10'b1010011001: angle = 16'b0001011101110111;
    10'b1010011010: angle = 16'b0001011101111110;
    10'b1010011011: angle = 16'b0001011110000101;
    10'b1010011100: angle = 16'b0001011110001100;
    10'b1010011101: angle = 16'b0001011110010100;
    10'b1010011110: angle = 16'b0001011110011011;
    10'b1010011111: angle = 16'b0001011110100010;
    10'b1010100000: angle = 16'b0001011110101001;
    10'b1010100001: angle = 16'b0001011110110000;
    10'b1010100010: angle = 16'b0001011110110111;
    10'b1010100011: angle = 16'b0001011110111110;
    10'b1010100100: angle = 16'b0001011111000101;
    10'b1010100101: angle = 16'b0001011111001101;
    10'b1010100110: angle = 16'b0001011111010100;
    10'b1010100111: angle = 16'b0001011111011011;
    10'b1010101000: angle = 16'b0001011111100010;
    10'b1010101001: angle = 16'b0001011111101001;
    10'b1010101010: angle = 16'b0001011111110000;
    10'b1010101011: angle = 16'b0001011111110111;
    10'b1010101100: angle = 16'b0001011111111110;
    10'b1010101101: angle = 16'b0001100000000101;
    10'b1010101110: angle = 16'b0001100000001100;
    10'b1010101111: angle = 16'b0001100000010011;
    10'b1010110000: angle = 16'b0001100000011010;
    10'b1010110001: angle = 16'b0001100000100001;
    10'b1010110010: angle = 16'b0001100000101000;
    10'b1010110011: angle = 16'b0001100000101111;
    10'b1010110100: angle = 16'b0001100000110110;
    10'b1010110101: angle = 16'b0001100000111101;
    10'b1010110110: angle = 16'b0001100001000100;
    10'b1010110111: angle = 16'b0001100001001011;
    10'b1010111000: angle = 16'b0001100001010010;
    10'b1010111001: angle = 16'b0001100001011001;
    10'b1010111010: angle = 16'b0001100001100000;
    10'b1010111011: angle = 16'b0001100001100111;
    10'b1010111100: angle = 16'b0001100001101110;
    10'b1010111101: angle = 16'b0001100001110101;
    10'b1010111110: angle = 16'b0001100001111100;
    10'b1010111111: angle = 16'b0001100010000011;
    10'b1011000000: angle = 16'b0001100010001010;
    10'b1011000001: angle = 16'b0001100010010000;
    10'b1011000010: angle = 16'b0001100010010111;
    10'b1011000011: angle = 16'b0001100010011110;
    10'b1011000100: angle = 16'b0001100010100101;
    10'b1011000101: angle = 16'b0001100010101100;
    10'b1011000110: angle = 16'b0001100010110011;
    10'b1011000111: angle = 16'b0001100010111010;
    10'b1011001000: angle = 16'b0001100011000001;
    10'b1011001001: angle = 16'b0001100011001000;
    10'b1011001010: angle = 16'b0001100011001110;
    10'b1011001011: angle = 16'b0001100011010101;
    10'b1011001100: angle = 16'b0001100011011100;
    10'b1011001101: angle = 16'b0001100011100011;
    10'b1011001110: angle = 16'b0001100011101010;
    10'b1011001111: angle = 16'b0001100011110001;
    10'b1011010000: angle = 16'b0001100011110111;
    10'b1011010001: angle = 16'b0001100011111110;
    10'b1011010010: angle = 16'b0001100100000101;
    10'b1011010011: angle = 16'b0001100100001100;
    10'b1011010100: angle = 16'b0001100100010011;
    10'b1011010101: angle = 16'b0001100100011001;
    10'b1011010110: angle = 16'b0001100100100000;
    10'b1011010111: angle = 16'b0001100100100111;
    10'b1011011000: angle = 16'b0001100100101110;
    10'b1011011001: angle = 16'b0001100100110101;
    10'b1011011010: angle = 16'b0001100100111011;
    10'b1011011011: angle = 16'b0001100101000010;
    10'b1011011100: angle = 16'b0001100101001001;
    10'b1011011101: angle = 16'b0001100101010000;
    10'b1011011110: angle = 16'b0001100101010110;
    10'b1011011111: angle = 16'b0001100101011101;
    10'b1011100000: angle = 16'b0001100101100100;
    10'b1011100001: angle = 16'b0001100101101010;
    10'b1011100010: angle = 16'b0001100101110001;
    10'b1011100011: angle = 16'b0001100101111000;
    10'b1011100100: angle = 16'b0001100101111111;
    10'b1011100101: angle = 16'b0001100110000101;
    10'b1011100110: angle = 16'b0001100110001100;
    10'b1011100111: angle = 16'b0001100110010011;
    10'b1011101000: angle = 16'b0001100110011001;
    10'b1011101001: angle = 16'b0001100110100000;
    10'b1011101010: angle = 16'b0001100110100111;
    10'b1011101011: angle = 16'b0001100110101101;
    10'b1011101100: angle = 16'b0001100110110100;
    10'b1011101101: angle = 16'b0001100110111010;
    10'b1011101110: angle = 16'b0001100111000001;
    10'b1011101111: angle = 16'b0001100111001000;
    10'b1011110000: angle = 16'b0001100111001110;
    10'b1011110001: angle = 16'b0001100111010101;
    10'b1011110010: angle = 16'b0001100111011100;
    10'b1011110011: angle = 16'b0001100111100010;
    10'b1011110100: angle = 16'b0001100111101001;
    10'b1011110101: angle = 16'b0001100111101111;
    10'b1011110110: angle = 16'b0001100111110110;
    10'b1011110111: angle = 16'b0001100111111101;
    10'b1011111000: angle = 16'b0001101000000011;
    10'b1011111001: angle = 16'b0001101000001010;
    10'b1011111010: angle = 16'b0001101000010000;
    10'b1011111011: angle = 16'b0001101000010111;
    10'b1011111100: angle = 16'b0001101000011101;
    10'b1011111101: angle = 16'b0001101000100100;
    10'b1011111110: angle = 16'b0001101000101010;
    10'b1011111111: angle = 16'b0001101000110001;
    10'b1100000000: angle = 16'b0001101000110111;
    10'b1100000001: angle = 16'b0001101000111110;
    10'b1100000010: angle = 16'b0001101001000100;
    10'b1100000011: angle = 16'b0001101001001011;
    10'b1100000100: angle = 16'b0001101001010001;
    10'b1100000101: angle = 16'b0001101001011000;
    10'b1100000110: angle = 16'b0001101001011110;
    10'b1100000111: angle = 16'b0001101001100101;
    10'b1100001000: angle = 16'b0001101001101011;
    10'b1100001001: angle = 16'b0001101001110010;
    10'b1100001010: angle = 16'b0001101001111000;
    10'b1100001011: angle = 16'b0001101001111111;
    10'b1100001100: angle = 16'b0001101010000101;
    10'b1100001101: angle = 16'b0001101010001100;
    10'b1100001110: angle = 16'b0001101010010010;
    10'b1100001111: angle = 16'b0001101010011001;
    10'b1100010000: angle = 16'b0001101010011111;
    10'b1100010001: angle = 16'b0001101010100101;
    10'b1100010010: angle = 16'b0001101010101100;
    10'b1100010011: angle = 16'b0001101010110010;
    10'b1100010100: angle = 16'b0001101010111001;
    10'b1100010101: angle = 16'b0001101010111111;
    10'b1100010110: angle = 16'b0001101011000101;
    10'b1100010111: angle = 16'b0001101011001100;
    10'b1100011000: angle = 16'b0001101011010010;
    10'b1100011001: angle = 16'b0001101011011001;
    10'b1100011010: angle = 16'b0001101011011111;
    10'b1100011011: angle = 16'b0001101011100101;
    10'b1100011100: angle = 16'b0001101011101100;
    10'b1100011101: angle = 16'b0001101011110010;
    10'b1100011110: angle = 16'b0001101011111000;
    10'b1100011111: angle = 16'b0001101011111111;
    10'b1100100000: angle = 16'b0001101100000101;
    10'b1100100001: angle = 16'b0001101100001011;
    10'b1100100010: angle = 16'b0001101100010010;
    10'b1100100011: angle = 16'b0001101100011000;
    10'b1100100100: angle = 16'b0001101100011110;
    10'b1100100101: angle = 16'b0001101100100101;
    10'b1100100110: angle = 16'b0001101100101011;
    10'b1100100111: angle = 16'b0001101100110001;
    10'b1100101000: angle = 16'b0001101100110111;
    10'b1100101001: angle = 16'b0001101100111110;
    10'b1100101010: angle = 16'b0001101101000100;
    10'b1100101011: angle = 16'b0001101101001010;
    10'b1100101100: angle = 16'b0001101101010000;
    10'b1100101101: angle = 16'b0001101101010111;
    10'b1100101110: angle = 16'b0001101101011101;
    10'b1100101111: angle = 16'b0001101101100011;
    10'b1100110000: angle = 16'b0001101101101001;
    10'b1100110001: angle = 16'b0001101101110000;
    10'b1100110010: angle = 16'b0001101101110110;
    10'b1100110011: angle = 16'b0001101101111100;
    10'b1100110100: angle = 16'b0001101110000010;
    10'b1100110101: angle = 16'b0001101110001000;
    10'b1100110110: angle = 16'b0001101110001111;
    10'b1100110111: angle = 16'b0001101110010101;
    10'b1100111000: angle = 16'b0001101110011011;
    10'b1100111001: angle = 16'b0001101110100001;
    10'b1100111010: angle = 16'b0001101110100111;
    10'b1100111011: angle = 16'b0001101110101110;
    10'b1100111100: angle = 16'b0001101110110100;
    10'b1100111101: angle = 16'b0001101110111010;
    10'b1100111110: angle = 16'b0001101111000000;
    10'b1100111111: angle = 16'b0001101111000110;
    10'b1101000000: angle = 16'b0001101111001100;
    10'b1101000001: angle = 16'b0001101111010010;
    10'b1101000010: angle = 16'b0001101111011001;
    10'b1101000011: angle = 16'b0001101111011111;
    10'b1101000100: angle = 16'b0001101111100101;
    10'b1101000101: angle = 16'b0001101111101011;
    10'b1101000110: angle = 16'b0001101111110001;
    10'b1101000111: angle = 16'b0001101111110111;
    10'b1101001000: angle = 16'b0001101111111101;
    10'b1101001001: angle = 16'b0001110000000011;
    10'b1101001010: angle = 16'b0001110000001001;
    10'b1101001011: angle = 16'b0001110000001111;
    10'b1101001100: angle = 16'b0001110000010110;
    10'b1101001101: angle = 16'b0001110000011100;
    10'b1101001110: angle = 16'b0001110000100010;
    10'b1101001111: angle = 16'b0001110000101000;
    10'b1101010000: angle = 16'b0001110000101110;
    10'b1101010001: angle = 16'b0001110000110100;
    10'b1101010010: angle = 16'b0001110000111010;
    10'b1101010011: angle = 16'b0001110001000000;
    10'b1101010100: angle = 16'b0001110001000110;
    10'b1101010101: angle = 16'b0001110001001100;
    10'b1101010110: angle = 16'b0001110001010010;
    10'b1101010111: angle = 16'b0001110001011000;
    10'b1101011000: angle = 16'b0001110001011110;
    10'b1101011001: angle = 16'b0001110001100100;
    10'b1101011010: angle = 16'b0001110001101010;
    10'b1101011011: angle = 16'b0001110001110000;
    10'b1101011100: angle = 16'b0001110001110110;
    10'b1101011101: angle = 16'b0001110001111100;
    10'b1101011110: angle = 16'b0001110010000010;
    10'b1101011111: angle = 16'b0001110010001000;
    10'b1101100000: angle = 16'b0001110010001110;
    10'b1101100001: angle = 16'b0001110010010100;
    10'b1101100010: angle = 16'b0001110010011010;
    10'b1101100011: angle = 16'b0001110010100000;
    10'b1101100100: angle = 16'b0001110010100101;
    10'b1101100101: angle = 16'b0001110010101011;
    10'b1101100110: angle = 16'b0001110010110001;
    10'b1101100111: angle = 16'b0001110010110111;
    10'b1101101000: angle = 16'b0001110010111101;
    10'b1101101001: angle = 16'b0001110011000011;
    10'b1101101010: angle = 16'b0001110011001001;
    10'b1101101011: angle = 16'b0001110011001111;
    10'b1101101100: angle = 16'b0001110011010101;
    10'b1101101101: angle = 16'b0001110011011011;
    10'b1101101110: angle = 16'b0001110011100000;
    10'b1101101111: angle = 16'b0001110011100110;
    10'b1101110000: angle = 16'b0001110011101100;
    10'b1101110001: angle = 16'b0001110011110010;
    10'b1101110010: angle = 16'b0001110011111000;
    10'b1101110011: angle = 16'b0001110011111110;
    10'b1101110100: angle = 16'b0001110100000100;
    10'b1101110101: angle = 16'b0001110100001001;
    10'b1101110110: angle = 16'b0001110100001111;
    10'b1101110111: angle = 16'b0001110100010101;
    10'b1101111000: angle = 16'b0001110100011011;
    10'b1101111001: angle = 16'b0001110100100001;
    10'b1101111010: angle = 16'b0001110100100110;
    10'b1101111011: angle = 16'b0001110100101100;
    10'b1101111100: angle = 16'b0001110100110010;
    10'b1101111101: angle = 16'b0001110100111000;
    10'b1101111110: angle = 16'b0001110100111110;
    10'b1101111111: angle = 16'b0001110101000011;
    10'b1110000000: angle = 16'b0001110101001001;
    10'b1110000001: angle = 16'b0001110101001111;
    10'b1110000010: angle = 16'b0001110101010101;
    10'b1110000011: angle = 16'b0001110101011010;
    10'b1110000100: angle = 16'b0001110101100000;
    10'b1110000101: angle = 16'b0001110101100110;
    10'b1110000110: angle = 16'b0001110101101100;
    10'b1110000111: angle = 16'b0001110101110001;
    10'b1110001000: angle = 16'b0001110101110111;
    10'b1110001001: angle = 16'b0001110101111101;
    10'b1110001010: angle = 16'b0001110110000011;
    10'b1110001011: angle = 16'b0001110110001000;
    10'b1110001100: angle = 16'b0001110110001110;
    10'b1110001101: angle = 16'b0001110110010100;
    10'b1110001110: angle = 16'b0001110110011001;
    10'b1110001111: angle = 16'b0001110110011111;
    10'b1110010000: angle = 16'b0001110110100101;
    10'b1110010001: angle = 16'b0001110110101010;
    10'b1110010010: angle = 16'b0001110110110000;
    10'b1110010011: angle = 16'b0001110110110110;
    10'b1110010100: angle = 16'b0001110110111011;
    10'b1110010101: angle = 16'b0001110111000001;
    10'b1110010110: angle = 16'b0001110111000111;
    10'b1110010111: angle = 16'b0001110111001100;
    10'b1110011000: angle = 16'b0001110111010010;
    10'b1110011001: angle = 16'b0001110111011000;
    10'b1110011010: angle = 16'b0001110111011101;
    10'b1110011011: angle = 16'b0001110111100011;
    10'b1110011100: angle = 16'b0001110111101001;
    10'b1110011101: angle = 16'b0001110111101110;
    10'b1110011110: angle = 16'b0001110111110100;
    10'b1110011111: angle = 16'b0001110111111001;
    10'b1110100000: angle = 16'b0001110111111111;
    10'b1110100001: angle = 16'b0001111000000101;
    10'b1110100010: angle = 16'b0001111000001010;
    10'b1110100011: angle = 16'b0001111000010000;
    10'b1110100100: angle = 16'b0001111000010101;
    10'b1110100101: angle = 16'b0001111000011011;
    10'b1110100110: angle = 16'b0001111000100000;
    10'b1110100111: angle = 16'b0001111000100110;
    10'b1110101000: angle = 16'b0001111000101100;
    10'b1110101001: angle = 16'b0001111000110001;
    10'b1110101010: angle = 16'b0001111000110111;
    10'b1110101011: angle = 16'b0001111000111100;
    10'b1110101100: angle = 16'b0001111001000010;
    10'b1110101101: angle = 16'b0001111001000111;
    10'b1110101110: angle = 16'b0001111001001101;
    10'b1110101111: angle = 16'b0001111001010010;
    10'b1110110000: angle = 16'b0001111001011000;
    10'b1110110001: angle = 16'b0001111001011101;
    10'b1110110010: angle = 16'b0001111001100011;
    10'b1110110011: angle = 16'b0001111001101000;
    10'b1110110100: angle = 16'b0001111001101110;
    10'b1110110101: angle = 16'b0001111001110011;
    10'b1110110110: angle = 16'b0001111001111001;
    10'b1110110111: angle = 16'b0001111001111110;
    10'b1110111000: angle = 16'b0001111010000100;
    10'b1110111001: angle = 16'b0001111010001001;
    10'b1110111010: angle = 16'b0001111010001111;
    10'b1110111011: angle = 16'b0001111010010100;
    10'b1110111100: angle = 16'b0001111010011001;
    10'b1110111101: angle = 16'b0001111010011111;
    10'b1110111110: angle = 16'b0001111010100100;
    10'b1110111111: angle = 16'b0001111010101010;
    10'b1111000000: angle = 16'b0001111010101111;
    10'b1111000001: angle = 16'b0001111010110101;
    10'b1111000010: angle = 16'b0001111010111010;
    10'b1111000011: angle = 16'b0001111010111111;
    10'b1111000100: angle = 16'b0001111011000101;
    10'b1111000101: angle = 16'b0001111011001010;
    10'b1111000110: angle = 16'b0001111011010000;
    10'b1111000111: angle = 16'b0001111011010101;
    10'b1111001000: angle = 16'b0001111011011010;
    10'b1111001001: angle = 16'b0001111011100000;
    10'b1111001010: angle = 16'b0001111011100101;
    10'b1111001011: angle = 16'b0001111011101010;
    10'b1111001100: angle = 16'b0001111011110000;
    10'b1111001101: angle = 16'b0001111011110101;
    10'b1111001110: angle = 16'b0001111011111011;
    10'b1111001111: angle = 16'b0001111100000000;
    10'b1111010000: angle = 16'b0001111100000101;
    10'b1111010001: angle = 16'b0001111100001011;
    10'b1111010010: angle = 16'b0001111100010000;
    10'b1111010011: angle = 16'b0001111100010101;
    10'b1111010100: angle = 16'b0001111100011011;
    10'b1111010101: angle = 16'b0001111100100000;
    10'b1111010110: angle = 16'b0001111100100101;
    10'b1111010111: angle = 16'b0001111100101010;
    10'b1111011000: angle = 16'b0001111100110000;
    10'b1111011001: angle = 16'b0001111100110101;
    10'b1111011010: angle = 16'b0001111100111010;
    10'b1111011011: angle = 16'b0001111101000000;
    10'b1111011100: angle = 16'b0001111101000101;
    10'b1111011101: angle = 16'b0001111101001010;
    10'b1111011110: angle = 16'b0001111101001111;
    10'b1111011111: angle = 16'b0001111101010101;
    10'b1111100000: angle = 16'b0001111101011010;
    10'b1111100001: angle = 16'b0001111101011111;
    10'b1111100010: angle = 16'b0001111101100100;
    10'b1111100011: angle = 16'b0001111101101010;
    10'b1111100100: angle = 16'b0001111101101111;
    10'b1111100101: angle = 16'b0001111101110100;
    10'b1111100110: angle = 16'b0001111101111001;
    10'b1111100111: angle = 16'b0001111101111111;
    10'b1111101000: angle = 16'b0001111110000100;
    10'b1111101001: angle = 16'b0001111110001001;
    10'b1111101010: angle = 16'b0001111110001110;
    10'b1111101011: angle = 16'b0001111110010011;
    10'b1111101100: angle = 16'b0001111110011001;
    10'b1111101101: angle = 16'b0001111110011110;
    10'b1111101110: angle = 16'b0001111110100011;
    10'b1111101111: angle = 16'b0001111110101000;
    10'b1111110000: angle = 16'b0001111110101101;
    10'b1111110001: angle = 16'b0001111110110011;
    10'b1111110010: angle = 16'b0001111110111000;
    10'b1111110011: angle = 16'b0001111110111101;
    10'b1111110100: angle = 16'b0001111111000010;
    10'b1111110101: angle = 16'b0001111111000111;
    10'b1111110110: angle = 16'b0001111111001100;
    10'b1111110111: angle = 16'b0001111111010001;
    10'b1111111000: angle = 16'b0001111111010111;
    10'b1111111001: angle = 16'b0001111111011100;
    10'b1111111010: angle = 16'b0001111111100001;
    10'b1111111011: angle = 16'b0001111111100110;
    10'b1111111100: angle = 16'b0001111111101011;
    10'b1111111101: angle = 16'b0001111111110000;
    10'b1111111110: angle = 16'b0001111111110101;
    10'b1111111111: angle = 16'b0001111111111010;
endcase
end
  
  
endmodule